entity empty is
end empty;